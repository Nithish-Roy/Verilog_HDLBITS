module top_module( input in, output out );
  assign out = ~(in); // out is assigned as not of in
endmodule
