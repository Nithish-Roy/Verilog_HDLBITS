module top_module( input in, output out );
assign out = in; // out is assigned to in which acts as a wire due to continous assignment
endmodule
