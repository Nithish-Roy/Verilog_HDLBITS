module top_module ( 
    input p1a, p1b, p1c, p1d, p1e, p1f,
    output p1y,
    input p2a, p2b, p2c, p2d,
    output p2y );
	  wire w1, w2, w3, w4;
    assign w1 = (p1a & p1b & p1c);
    assign w2 = (p1d & p1e & p1f);
    assign p1y = (w1 | w2);
    assign w3 = (p2a & p2b);
    assign w4 = (p2c & p2d);
    assign p2y = (w3 | w4);

endmodule
/* the code was written based on the image : https://hdlbits.01xz.net/mw/images/e/e1/7458.png*/
