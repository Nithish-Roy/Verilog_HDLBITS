module top_module(
    output zero
);// Module body starts after semicolon
assign zero = 1'b0;    // zero is assigned to 0
endmodule
